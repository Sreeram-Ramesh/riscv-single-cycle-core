`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Designer: Sreeram R 
// 
// Create Date: 08/16/2025 05:58:40 PM
// Design Name: Vanilla RV32I
// Module Name: riscv32i_cpu
// Project Name: 
// Target Devices: Zynq 7000
// Tool Versions: 
// Description: 
// 
// Dependencies: A hex file with instructions to be loaded into the instruction
//               memory.
// 
// Revision: v01
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module riscv32i_cpu (
    input         clk, reset,
    input         Stall,
    input         Ext_MemWrite,
    input  [31:0] Ext_WriteData, Ext_DataAdr,
    output        MemWrite,
    output [31:0] WriteData, DataAdr, ReadData,
    output [31:0] PC, Result
);

wire [31:0] Instr;
wire [31:0] DataAdr_rv32, WriteData_rv32;
wire        MemWrite_rv32;

// instantiate processor and memories
riscv_cpu rvcpu    (clk, reset, Stall, PC, Instr,
                    MemWrite_rv32, DataAdr_rv32,
                    WriteData_rv32, ReadData, Result);
instr_mem instrmem (PC, Instr);
data_mem  datamem  (clk, MemWrite, Stall, Instr[14:12], DataAdr, WriteData, ReadData);

assign MemWrite  = (Ext_MemWrite && reset) ? 1 : MemWrite_rv32;
assign WriteData = (Ext_MemWrite && reset) ? Ext_WriteData : WriteData_rv32;
assign DataAdr   = reset ? Ext_DataAdr : DataAdr_rv32;

endmodule
